.title KiCad test

.include ./inverter.ngcir

* Adding the source
a1 [I_BUS] input_vector
.model input_vector d_source(input_file = "testdata.txt")

* Then convert this to analog
adac0 [I_BUS ] [ A ] dac
.model dac dac_bridge(out_low = 0 out_high = 1 out_undef = 0.5 input_load = 5.0e-12 t_rise = 0.11e-9 t_fall = 0.1e-9)


Vvss vss 0 0

Xinv A Z inverter
.tran 1e-5 10e-9
.control
set wr_singlescale
set wr_vecnames
run
wrdata inverter_A.csv v(A)
wrdata inverter_Z.csv v(Z)
.endc

.end
